module triStateBuffer(
		input a , c ,
		output f
	);

	bufif1(f , a , c);
endmodule
